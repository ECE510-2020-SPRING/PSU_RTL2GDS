module MUX21X2 ( input A1, input A2, input S0, output Y );
   MUX21X2_HVT mux21x2_inst (.A1(A1), .A2(A2), .S0(S0), .Y(Y) );
endmodule

