// A simple AND gate

module simple_and (ain, bin, cout );

input ain, bin ;

output cout;

assign cout = ain & bin;

endmodule
